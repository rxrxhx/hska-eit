/* Verilog model created from schematic test.sch -- Sep 20, 2018 00:31 */

module test( O );
output O;



defparam I1.NOM_FREQ="2.08";
OSCH I1 ( .OSC(O) );

endmodule // test
